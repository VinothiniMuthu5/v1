module test();
  initial begin
    display("Hello");
  end
endmodule
